magic
tech scmos
timestamp 1569736965
<< nwell >>
rect -19 -13 9 11
<< polysilicon >>
rect -6 3 -4 6
rect -6 -2 -4 0
<< pdiffusion >>
rect -7 0 -6 3
rect -4 0 -3 3
<< metal1 >>
rect -2 6 8 9
rect -11 -3 -8 -1
rect -18 -6 -8 -3
rect -2 -8 1 -1
rect -9 -12 -2 -9
<< ptransistor >>
rect -6 0 -4 3
<< polycontact >>
rect -6 6 -2 10
<< pdcontact >>
rect -11 -1 -7 3
rect -3 -1 1 3
<< nsubstratencontact >>
rect -2 -12 2 -8
<< labels >>
rlabel metal1 -8 -11 -8 -11 1 VDD
rlabel metal1 -17 -5 -17 -5 3 GND
rlabel metal1 6 7 6 7 6 GATE
<< end >>
