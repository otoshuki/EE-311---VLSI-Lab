Question 6 - 8-Bit Register
*Guining Pertin - 170102027

*Default parameters
.MODEL PMOS1 PMOS
.MODEL NMOS1 NMOS

*CMOS NOT Gate
.SUBCKT NOT VDD GND IN OUT
M1 OUT IN GND GND NMOS1
M2 OUT IN VDD VDD PMOS1
.ENDS NOT

*CMOS 2-Input NAND Gate
.SUBCKT NAND2 VDD GND A B OUT
M1 OUT A 1 1 NMOS1
M2 1 B GND GND NMOS1
M3 OUT A VDD VDD PMOS1
M4 OUT B VDD VDD PMOS1
.ENDS NAND

*CMOS 3-Input NAND Gate
.SUBCKT NAND3 VDD GND A B C OUT
M1 OUT A 1 1 NMOS1
M2 1 B 2 2 NMOS1
M3 2 C GND GND NMOS1
M4 OUT A VDD VDD PMOS1
M5 OUT B VDD VDD PMOS1
M6 OUT C VDD VDD PMOS1
.ENDS NAND3

*Positive Edge Triggered D Flip Flop
.SUBCKT DFLIP VDD GND CLK D Q
X1 VDD GND N4 N2 N1 NAND2
X2 VDD GND N1 CLK N2 NAND2
X3 VDD GND N2 CLK N4 N3 NAND3
X4 VDD GND N3 D N4 NAND2
X5 VDD GND N2 QP Q NAND2
X6 VDD GND N3 Q QP NAND2
.ENDS DFLIP

*8-Bit Register
VD VDD GND DC 5
X0 VDD GND CLK D0 Q0 DFLIP
X1 VDD GND CLK D1 Q1 DFLIP
X2 VDD GND CLK D2 Q2 DFLIP
X3 VDD GND CLK D3 Q3 DFLIP
X4 VDD GND CLK D4 Q4 DFLIP
X5 VDD GND CLK D5 Q5 DFLIP
X6 VDD GND CLK D6 Q6 DFLIP
X7 VDD GND CLK D7 Q7 DFLIP

*Clock
VCLK CLK GND DC 0 AC 0 PULSE(0 4 1.2 0.2 0.2 1 1)

*Input to store
V0 D0 GND DC 0 AC 0 PULSE(0 5 5 0 0 5 5)
V1 D1 GND DC 0 AC 0 PULSE(5 0 5 0 0 5 5)
V2 D2 GND DC 0 AC 0 PULSE(0 5 5 0 0 5 5)
V3 D3 GND DC 0 AC 0 PULSE(5 0 5 0 0 5 5)
V4 D4 GND DC 0 AC 0 PULSE(0 5 5 0 0 5 5)
V5 D5 GND DC 0 AC 0 PULSE(0 5 5 0 0 5 5)
V6 D6 GND DC 0 AC 0 PULSE(0 5 5 0 0 5 5)
V7 D7 GND DC 0 AC 0 PULSE(5 0 5 0 0 5 5)

.control

tran 10m 10 2
plot D0 
plot D1 

.endc

.end
