Question 5 - 2-Input CMOS XOR Gate
*Guining Pertin - 170102027

*Default parameters
.MODEL PMOS1 PMOS
.MODEL NMOS1 NMOS

*CMOS NOT Gate
.SUBCKT NOT VDD GND IN OUT
M1 OUT IN GND GND NMOS1
M2 OUT IN VDD VDD PMOS1
C1 OUT GND 0.1u
.ENDS NOT

*CMOS NAND Gate
.SUBCKT NAND VDD GND A B OUT
M1 OUT A 1 1 NMOS1
M2 1 B GND GND NMOS1
M3 OUT A VDD VDD PMOS1
M4 OUT B VDD VDD PMOS1
.ENDS NAND

*CMOS XOR Gate
V1 VDD GND DC 5
X1 VDD GND A AP NOT
X2 VDD GND B BP NOT
X3 VDD GND AP B N1 NAND
X4 VDD GND A BP N2 NAND
X5 VDD GND N1 N2 OUT NAND

*Pulse inputs for each ABC combination
VA A GND DC 0 AC 0 PULSE(0 5 2 0 0 2 4)
VB B GND DC 0 AC 0 PULSE(0 5 1 0 0 1 2)

.control

tran 10m 4
plot OUT ylabel 'Output(0110)'

.endc

.end
