* SPICE3 file created from q5_nand.ext - technology: scmos
*Question 5 - 3-input NAND
*Guining Pertin - 170102027

.option scale=1u
.MODEL nfet NMOS
.MODEL pfet PMOS

*MAGIC extractions
*PMOS
M1000 OUT A VDD VDD pfet w=3 l=2 ad=41 pd=38 as=41 ps=38
M1001 OUT B VDD VDD pfet w=3 l=2 ad=0 pd=0 as=0 ps=0
M1002 OUT C VDD VDD pfet w=3 l=2 ad=0 pd=0 as=0 ps=0
*NMOS
M1003 OUT A inter1 GND nfet w=3 l=2 ad=18 pd=18 as=19 ps=18
M1004 inter1 B inter2 GND nfet w=3 l=2 ad=18 pd=18 as=0 ps=0
M1005 inter2 C GND GND nfet w=3 l=2 ad=19 pd=18 as=0 ps=0
*Parasitics
C0 OUT VDD 7.7fF
C1 VDD GND 8.1fF

*Voltage Sources
VD VDD GND DC 5
VA A GND DC 0 AC 0 PULSE(0 5 3.8 0.2 0.2 3.8 8)
VB B GND DC 0 AC 0 PULSE(0 5 1.8 0.2 0.2 1.8 4)
VC C GND DC 0 AC 0 PULSE(0 5 0.8 0.2 0.2 0.8 2)

.CONTROL

TRAN 10m 8
PLOT C OUT ylabel 'LSB/OUTPUT'

.ENDC

.END
