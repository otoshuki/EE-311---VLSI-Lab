magic
tech scmos
timestamp 1569753433
<< nwell >>
rect -11 6 19 37
<< polysilicon >>
rect -5 14 -3 16
rect 3 14 5 16
rect 11 14 13 16
rect -5 8 -3 11
rect 3 8 5 11
rect 11 8 13 11
rect -5 4 -4 8
rect 3 4 4 8
rect 11 4 12 8
rect -5 1 -3 4
rect 3 1 5 4
rect 11 1 13 4
rect -5 -4 -3 -2
rect 3 -4 5 -2
rect 11 -4 13 -2
<< ndiffusion >>
rect -6 -2 -5 1
rect -3 -2 3 1
rect 5 -2 11 1
rect 13 -2 14 1
<< pdiffusion >>
rect -6 11 -5 14
rect -3 11 -2 14
rect 2 11 3 14
rect 5 11 6 14
rect 10 11 11 14
rect 13 11 14 14
<< metal1 >>
rect -11 31 -10 35
rect -6 31 -2 35
rect 2 31 7 35
rect 11 31 19 35
rect -10 25 10 28
rect -10 15 -7 25
rect -1 15 2 18
rect 7 15 10 25
rect 15 15 18 18
rect -10 7 -7 11
rect -18 4 -7 7
rect 0 4 1 8
rect 8 4 9 8
rect 16 4 17 8
rect -10 1 -7 4
rect 15 -7 18 -3
rect -11 -11 -10 -7
rect -6 -11 -2 -7
rect 2 -11 6 -7
rect 10 -11 14 -7
rect 18 -11 19 -7
<< metal2 >>
rect 11 31 19 35
rect 7 21 10 31
rect 2 18 14 21
<< ntransistor >>
rect -5 -2 -3 1
rect 3 -2 5 1
rect 11 -2 13 1
<< ptransistor >>
rect -5 11 -3 14
rect 3 11 5 14
rect 11 11 13 14
<< polycontact >>
rect -4 4 0 8
rect 4 4 8 8
rect 12 4 16 8
<< ndcontact >>
rect -10 -3 -6 1
rect 14 -3 18 1
<< pdcontact >>
rect -10 11 -6 15
rect -2 11 2 15
rect 6 11 10 15
rect 14 11 18 15
<< m2contact >>
rect 7 31 11 35
rect -2 18 2 22
rect 14 18 18 22
<< psubstratepcontact >>
rect -10 -11 -6 -7
rect -2 -11 2 -7
rect 6 -11 10 -7
rect 14 -11 18 -7
<< nsubstratencontact >>
rect -10 31 -6 35
rect -2 31 2 35
<< labels >>
rlabel polycontact 0 6 0 6 1 A
rlabel polycontact 8 6 8 6 1 B
rlabel polycontact 16 6 16 6 7 C
rlabel metal1 5 -9 5 -9 1 GND
rlabel metal1 -16 5 -16 5 3 OUT
rlabel metal2 16 33 16 33 6 VDD
rlabel ndiffusion 0 -1 0 -1 1 inter1
rlabel ndiffusion 8 -1 8 -1 1 inter2
<< end >>
