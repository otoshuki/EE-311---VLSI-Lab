Question 6 - 16-Bit Counter
*Guining Pertin - 170102027

*Default parameters
.MODEL PMOS1 PMOS
.MODEL NMOS1 NMOS

*CMOS NOT Gate
.SUBCKT NOT VDD GND IN OUT
M1 OUT IN GND GND NMOS1
M2 OUT IN VDD VDD PMOS1
.ENDS NOT

*CMOS 3-Input NAND Gate
.SUBCKT NAND3 VDD GND A B C OUT
M1 OUT A 1 1 NMOS1
M2 1 B 2 2 NMOS1
M3 2 C GND GND NMOS1
M4 OUT A VDD VDD PMOS1
M5 OUT B VDD VDD PMOS1
M6 OUT C VDD VDD PMOS1
.ENDS NAND3

*Positive Edge Triggered D Flip Flop
.SUBCKT DFLIP VDD GND CLK D Q QP PRESET CLEAR
X1 VDD GND N4 N2 PRESET N1 NAND3
X2 VDD GND N1 CLK CLEAR N2 NAND3
X3 VDD GND N2 CLK N4 N3 NAND3
X4 VDD GND N3 D CLEAR N4 NAND3
X5 VDD GND N2 QP PRESET Q NAND3
X6 VDD GND N3 Q CLEAR QP NAND3
.ENDS DFLIP

*16-Bit Binary Ripple Counter
VD VDD GND DC 5
X0 VDD GND CLK QP0 Q0 QP0 PRESET CLEAR DFLIP
X1 VDD GND QP0 QP1 Q1 QP1 PRESET CLEAR DFLIP
X2 VDD GND QP1 QP2 Q2 QP2 PRESET CLEAR DFLIP
X3 VDD GND QP2 QP3 Q3 QP3 PRESET CLEAR DFLIP
X4 VDD GND QP3 QP4 Q4 QP4 PRESET CLEAR DFLIP
X5 VDD GND QP4 QP5 Q5 QP5 PRESET CLEAR DFLIP
X6 VDD GND QP5 QP6 Q6 QP6 PRESET CLEAR DFLIP
X7 VDD GND QP6 QP7 Q7 QP7 PRESET CLEAR DFLIP
X8 VDD GND QP7 QP8 Q8 QP8 PRESET CLEAR DFLIP
X9 VDD GND QP8 QP9 Q9 QP9 PRESET CLEAR DFLIP
X10 VDD GND QP9 QP10 Q10 QP10 PRESET CLEAR DFLIP
X11 VDD GND QP10 QP11 Q11 QP11 PRESET CLEAR DFLIP
X12 VDD GND QP11 QP12 Q12 QP12 PRESET CLEAR DFLIP
X13 VDD GND QP12 QP13 Q13 QP13 PRESET CLEAR DFLIP
X14 VDD GND QP13 QP14 Q14 QP14 PRESET CLEAR DFLIP
X15 VDD GND QP14 QP15 Q15 QP15 PRESET CLEAR DFLIP
X16 VDD GND QP15 QP16 Q16 QP16 PRESET CLEAR DFLIP
X17 VDD GND QP16 QP17 Q17 QP17 PRESET CLEAR DFLIP

*Clock
VCLK CLK GND DC 0 AC 0 PULSE(0 4 1 0 0 1 2)
VPRE PRESET GND DC 5
VCLE CLEAR  GND DC 5

*Preset
.control

tran 10m 10
plot CLK
print all

.endc

.end
