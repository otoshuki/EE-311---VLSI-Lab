magic
tech scmos
timestamp 1569738269
<< nwell >>
rect -13 3 7 19
<< polysilicon >>
rect -5 8 -3 10
rect -5 2 -3 5
rect -4 -2 -3 2
rect -5 -5 -3 -2
rect -5 -10 -3 -8
<< ndiffusion >>
rect -6 -8 -5 -5
rect -3 -8 -2 -5
<< pdiffusion >>
rect -6 5 -5 8
rect -3 5 -2 8
<< metal1 >>
rect -12 14 -10 18
rect -6 14 -2 18
rect 2 14 6 18
rect -10 9 -7 14
rect -1 2 2 5
rect -13 -2 -8 2
rect -1 -2 7 2
rect -1 -5 2 -2
rect -10 -14 -7 -9
rect -12 -18 -10 -14
rect -6 -18 -2 -14
rect 2 -18 6 -14
<< ntransistor >>
rect -5 -8 -3 -5
<< ptransistor >>
rect -5 5 -3 8
<< polycontact >>
rect -8 -2 -4 2
<< ndcontact >>
rect -10 -9 -6 -5
rect -2 -9 2 -5
<< pdcontact >>
rect -10 5 -6 9
rect -2 5 2 9
<< psubstratepcontact >>
rect -10 -18 -6 -14
rect -2 -18 2 -14
<< nsubstratencontact >>
rect -10 14 -6 18
rect -2 14 2 18
<< labels >>
rlabel metal1 -12 0 -12 0 3 A
rlabel metal1 6 0 6 0 7 A_BAR
rlabel metal1 4 16 4 16 6 VDD
rlabel metal1 4 -16 4 -16 8 GND
<< end >>
