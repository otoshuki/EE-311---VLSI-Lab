magic
tech scmos
timestamp 1569754665
<< nwell >>
rect -9 3 21 21
<< polysilicon >>
rect -3 11 -1 13
rect 5 11 7 13
rect 13 11 15 13
rect -3 5 -1 8
rect 5 5 7 8
rect 13 5 15 8
rect -3 1 -2 5
rect 5 1 6 5
rect 13 1 14 5
rect -3 -2 -1 1
rect 5 -2 7 1
rect 13 -2 15 1
rect -3 -7 -1 -5
rect 5 -7 7 -5
rect 13 -7 15 -5
<< ndiffusion >>
rect -4 -5 -3 -2
rect -1 -5 0 -2
rect 4 -5 5 -2
rect 7 -5 8 -2
rect 12 -5 13 -2
rect 15 -5 16 -2
<< pdiffusion >>
rect -4 8 -3 11
rect -1 8 5 11
rect 7 8 13 11
rect 15 8 16 11
<< metal1 >>
rect -9 16 -8 20
rect -4 16 0 20
rect 4 16 8 20
rect 12 16 16 20
rect 20 16 21 20
rect 17 12 20 16
rect -8 5 -5 8
rect -17 1 -5 5
rect 2 1 3 5
rect 10 1 11 5
rect 18 1 19 5
rect -8 -2 -5 1
rect -8 -15 -5 -6
rect 1 -8 4 -6
rect 9 -15 12 -6
rect 17 -8 20 -6
rect -8 -18 12 -15
rect -9 -25 -8 -21
rect -4 -25 0 -21
rect 4 -25 9 -21
<< metal2 >>
rect 5 -12 17 -9
rect 9 -21 12 -12
rect 13 -25 22 -21
<< ntransistor >>
rect -3 -5 -1 -2
rect 5 -5 7 -2
rect 13 -5 15 -2
<< ptransistor >>
rect -3 8 -1 11
rect 5 8 7 11
rect 13 8 15 11
<< polycontact >>
rect -2 1 2 5
rect 6 1 10 5
rect 14 1 18 5
<< ndcontact >>
rect -8 -6 -4 -2
rect 0 -6 4 -2
rect 8 -6 12 -2
rect 16 -6 20 -2
<< pdcontact >>
rect -8 8 -4 12
rect 16 8 20 12
<< m2contact >>
rect 1 -12 5 -8
rect 17 -12 21 -8
rect 9 -25 13 -21
<< psubstratepcontact >>
rect -8 -25 -4 -21
rect 0 -25 4 -21
<< nsubstratencontact >>
rect -8 16 -4 20
rect 0 16 4 20
rect 8 16 12 20
rect 16 16 20 20
<< labels >>
rlabel metal2 17 -23 17 -23 8 GND
rlabel polycontact 2 2 2 2 1 A
rlabel polycontact 10 2 10 2 1 B
rlabel polycontact 18 3 18 3 7 C
rlabel metal1 14 18 14 18 5 VDD
rlabel pdiffusion 2 9 2 9 1 inter1
rlabel pdiffusion 10 9 10 9 1 inter2
rlabel metal1 -12 2 -12 2 3 OUT
<< end >>
