Question 10 - Two Stage Differential Amplifier
*Guining Pertin - 170102027

*Default parameters
.MODEL PMOS1 PMOS
.MODEL NMOS1 NMOS

*Single Stage Amplifier
.SUBCKT AMP VDD GND VIN1 VIN2 D5 D6
M0 D0 VB1 VDD VDD PMOS1
M1 D1 VIN1 D0 D0 PMOS1
M2 D2 VIN2 D0 D0 PMOS1
M3 D1 VB2 GND GND NMOS1
M4 D2 VB2 GND GND NMOS1
M5 D5 VB3 D1 D1 NMOS1
M6 D6 VB3 D2 D2 NMOS1
M7 D5 VB4 S7 S7 PMOS1
M8 D6 VB4 S8 S8 PMOS1
M9 S7 VB5 VDD VDD PMOS1
M10 S8 VB5 VDD VDD PMOS1
*Bias Voltages
V1 VB1 GND DC 3
V2 VB2 GND DC 3
V3 VB3 GND DC 3
V4 VB4 GND DC 3
V5 VB5 GND DC 3
.ENDS AMP

*Two Stage Amplifier
VD VDD GND DC 5
VIN VIN1 VIN2 DC 3 AC 3 SIN(0 30m 40k 0 0)
X1 VDD GND VIN1 VIN2 OUT1 OUT2 AMP
X2 VDD GND OUT1 OUT2 OUT3 OUT4 AMP

.control

op
tran 10u 10m
display
print all
*plot V(D5)

.endc

.end
