magic
tech scmos
timestamp 1569760954
<< nwell >>
rect -14 6 88 34
<< polysilicon >>
rect -8 13 -6 15
rect 8 13 10 15
rect 16 13 18 15
rect 32 13 34 15
rect 40 13 42 15
rect 56 13 58 15
rect 64 13 66 15
rect 80 13 82 16
rect -8 7 -6 10
rect 8 7 10 10
rect 16 7 18 10
rect 32 7 34 10
rect -7 3 -6 7
rect 9 3 10 7
rect 17 3 18 7
rect 33 3 34 7
rect -8 0 -6 3
rect 8 0 10 3
rect 16 0 18 3
rect 32 0 34 3
rect 40 7 42 10
rect 56 7 58 10
rect 64 7 66 10
rect 80 7 82 10
rect 40 3 41 7
rect 56 3 57 7
rect 64 3 65 7
rect 80 3 81 7
rect 40 0 42 3
rect 56 0 58 3
rect 64 0 66 3
rect 80 0 82 3
rect -8 -5 -6 -3
rect 8 -5 10 -3
rect 16 -5 18 -3
rect 32 -5 34 -3
rect 40 -5 42 -3
rect 56 -5 58 -3
rect 64 -5 66 -3
rect 80 -5 82 -3
<< ndiffusion >>
rect -9 -3 -8 0
rect -6 -3 -5 0
rect 7 -3 8 0
rect 10 -3 16 0
rect 18 -3 19 0
rect 31 -3 32 0
rect 34 -3 40 0
rect 42 -3 43 0
rect 55 -3 56 0
rect 58 -3 64 0
rect 66 -3 67 0
rect 79 -3 80 0
rect 82 -3 83 0
<< pdiffusion >>
rect -9 10 -8 13
rect -6 10 -5 13
rect 7 10 8 13
rect 10 10 11 13
rect 15 10 16 13
rect 18 10 19 13
rect 31 10 32 13
rect 34 10 35 13
rect 39 10 40 13
rect 42 10 43 13
rect 55 10 56 13
rect 58 10 59 13
rect 63 10 64 13
rect 66 10 67 13
rect 79 10 80 13
rect 82 10 83 13
<< metal1 >>
rect -9 29 -5 33
rect 79 29 83 33
rect -13 23 -9 29
rect -13 14 -9 19
rect 3 24 23 27
rect 3 14 6 24
rect 11 14 14 17
rect 20 14 23 24
rect 27 25 47 27
rect 27 24 43 25
rect 27 14 30 24
rect 35 14 39 17
rect 44 14 47 21
rect 51 24 71 27
rect 51 14 54 24
rect 60 14 63 17
rect 68 14 71 24
rect 83 23 87 29
rect 83 14 87 19
rect -4 7 -1 10
rect 20 7 23 10
rect 51 7 54 10
rect 75 7 78 10
rect -22 3 -11 7
rect -4 3 5 7
rect 20 3 29 7
rect 45 3 54 7
rect 69 3 78 7
rect 85 3 96 7
rect -19 -7 -16 3
rect -4 0 -1 3
rect -12 -7 -9 -4
rect 3 -7 6 -4
rect -12 -11 6 -7
rect -1 -20 3 -11
rect 13 -14 16 3
rect 20 0 23 3
rect 51 0 54 3
rect 27 -7 30 -4
rect 44 -7 47 -4
rect 58 -7 61 3
rect 75 0 78 3
rect 68 -11 71 -4
rect 83 -7 87 -4
rect 75 -11 87 -7
rect 90 -14 93 3
rect 13 -17 93 -14
rect -9 -24 15 -20
rect 19 -24 42 -20
rect 46 -24 59 -20
rect 63 -24 71 -20
<< metal2 >>
rect -1 29 75 33
rect 11 21 15 29
rect 35 21 39 29
rect 44 14 47 21
rect 59 21 63 29
rect 43 10 47 14
rect 44 -7 47 10
rect 10 -11 27 -7
rect 47 -11 52 -7
rect -19 -15 -16 -11
rect 58 -15 61 -11
rect -19 -18 61 -15
rect 71 -20 75 -11
rect 75 -24 86 -20
<< ntransistor >>
rect -8 -3 -6 0
rect 8 -3 10 0
rect 16 -3 18 0
rect 32 -3 34 0
rect 40 -3 42 0
rect 56 -3 58 0
rect 64 -3 66 0
rect 80 -3 82 0
<< ptransistor >>
rect -8 10 -6 13
rect 8 10 10 13
rect 16 10 18 13
rect 32 10 34 13
rect 40 10 42 13
rect 56 10 58 13
rect 64 10 66 13
rect 80 10 82 13
<< polycontact >>
rect -11 3 -7 7
rect 5 3 9 7
rect 13 3 17 7
rect 29 3 33 7
rect 41 3 45 7
rect 57 3 61 7
rect 65 3 69 7
rect 81 3 85 7
<< ndcontact >>
rect -13 -4 -9 0
rect -5 -4 -1 0
rect 3 -4 7 0
rect 19 -4 23 0
rect 27 -4 31 0
rect 43 -4 47 0
rect 51 -4 55 0
rect 67 -4 71 0
rect 75 -4 79 0
rect 83 -4 87 0
<< pdcontact >>
rect -13 10 -9 14
rect -5 10 -1 14
rect 3 10 7 14
rect 11 10 15 14
rect 19 10 23 14
rect 27 10 31 14
rect 35 10 39 14
rect 43 10 47 14
rect 51 10 55 14
rect 59 10 63 14
rect 67 10 71 14
rect 75 10 79 14
rect 83 10 87 14
<< m2contact >>
rect -5 29 -1 33
rect 75 29 79 33
rect 11 17 15 21
rect 43 21 47 25
rect 35 17 39 21
rect 59 17 63 21
rect -19 -11 -15 -7
rect 6 -11 10 -7
rect 27 -11 31 -7
rect 43 -11 47 -7
rect 58 -11 62 -7
rect 71 -11 75 -7
rect 71 -24 75 -20
<< psubstratepcontact >>
rect -13 -24 -9 -20
rect 15 -24 19 -20
rect 42 -24 46 -20
rect 59 -24 63 -20
<< nsubstratencontact >>
rect -13 29 -9 33
rect 83 29 87 33
rect -13 19 -9 23
rect 83 19 87 23
<< labels >>
rlabel metal1 74 5 74 5 1 B_BAR
rlabel metal1 -20 5 -20 5 3 A
rlabel metal1 94 5 94 5 7 B
rlabel metal1 24 5 24 5 1 N1
rlabel metal2 50 -9 50 -9 1 OUT
rlabel metal2 81 -22 81 -22 1 GND
rlabel ndiffusion 12 -2 12 -2 1 inter1
rlabel ndiffusion 62 -1 62 -1 1 inter2
rlabel ndiffusion 37 -2 37 -2 1 inter3
rlabel metal1 49 5 49 5 1 N2
rlabel metal1 2 5 2 5 1 A_BAR
rlabel metal2 37 31 37 31 1 VDD
<< end >>
