magic
tech scmos
timestamp 1569761636
<< polysilicon >>
rect 0 3 2 6
rect 0 -2 2 0
<< ndiffusion >>
rect -1 0 0 3
rect 2 0 3 3
<< metal1 >>
rect -7 6 -1 10
rect -5 -6 -2 -1
rect 4 -5 7 -1
rect 8 -9 12 -5
<< ntransistor >>
rect 0 0 2 3
<< polycontact >>
rect -1 6 3 10
<< ndcontact >>
rect -5 -1 -1 3
rect 3 -1 7 3
<< psubstratepcontact >>
rect 4 -9 8 -5
<< labels >>
rlabel metal1 -5 8 -5 8 4 GATE
rlabel metal1 -3 -4 -3 -4 2 VDD
rlabel metal1 9 -7 9 -7 8 GND
<< end >>
