Question 6 - 16-Bit Counter
*Guining Pertin - 170102027

*Default parameters
.MODEL PMOS1 PMOS
.MODEL NMOS1 NMOS

*CMOS NOT Gate
.SUBCKT NOT VDD GND IN OUT
M1 OUT IN GND GND NMOS1
M2 OUT IN VDD VDD PMOS1
.ENDS NOT

*CMOS 2-Input NAND Gate
.SUBCKT NAND2 VDD GND A B OUT
M1 OUT A 1 1 NMOS1
M2 1 B GND GND NMOS1
M3 OUT A VDD VDD PMOS1
M4 OUT B VDD VDD PMOS1
.ENDS NAND

*CMOS 3-Input NAND Gate
.SUBCKT NAND3 VDD GND A B C OUT
M1 OUT A 1 1 NMOS1
M2 1 B 2 2 NMOS1
M3 2 C GND GND NMOS1
M4 OUT A VDD VDD PMOS1
M5 OUT B VDD VDD PMOS1
M6 OUT C VDD VDD PMOS1
.ENDS NAND3

*Positive Edge Triggered D Flip Flop
.SUBCKT DFLIP VDD GND CLK D Q QP PRESET
X1 VDD GND N4 N2 PRESET N1 NAND3
X2 VDD GND N1 CLK N2 NAND2
X3 VDD GND N2 CLK N4 N3 NAND3
X4 VDD GND N3 D N4 NAND2
X5 VDD GND N2 QP PRESET Q NAND3
X6 VDD GND N3 Q QP NAND2
.ENDS DFLIP

*3-Bit Binary Ripple Counter
VD VDD GND DC 5
X0 VDD GND CLK QP0 Q0 QP0 PRESET DFLIP
X1 VDD GND QP0 QP1 Q1 QP1 PRESET DFLIP
X2 VDD GND QP1 QP2 Q2 QP2 PRESET DFLIP

*Clock
VCLK CLK GND DC 0 AC 0 PULSE(0 5 1 0 0 1 2)
VPRE PRESET GND DC 0 AC 0 PULSE(0 5 0.5 0 0 10 10)

*Preset
.control

tran 10m 10
plot Q0 Q1

.endc

.end
